
module button (
	buttons_write,
	clk_clk,
	reset_reset_n);	

	input	[7:0]	buttons_write;
	input		clk_clk;
	input		reset_reset_n;
endmodule
