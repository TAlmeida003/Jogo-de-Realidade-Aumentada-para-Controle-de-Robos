// Arquitetura.v

// Generated using ACDS version 23.1 993

`timescale 1 ps / 1 ps
module Arquitetura (
		input  wire        a_button_export,           //           a_button.export
		input  wire        b_button_export,           //           b_button.export
		input  wire        clk_clk,                   //                clk.clk
		output wire [31:0] data_a_export,             //             data_a.export
		output wire [31:0] data_b_export,             //             data_b.export
		input  wire [3:0]  direction_analogic_export, // direction_analogic.export
		input  wire        reset_reset_n,             //              reset.reset_n
		output wire        reset_pulsecounter_export, // reset_pulsecounter.export
		input  wire        screen_export,             //             screen.export
		input  wire        select_button_export,      //      select_button.export
		input  wire        start_button_export,       //       start_button.export
		input  wire        tl_button_export,          //          tl_button.export
		input  wire        tr_button_export,          //          tr_button.export
		input  wire        wrfull_export,             //             wrfull.export
		output wire        wrreg_export,              //              wrreg.export
		input  wire        x_button_export,           //           x_button.export
		input  wire        y_button_export            //           y_button.export
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [16:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [16:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_data_a_s1_chipselect;                      // mm_interconnect_0:data_A_s1_chipselect -> data_A:chipselect
	wire  [31:0] mm_interconnect_0_data_a_s1_readdata;                        // data_A:readdata -> mm_interconnect_0:data_A_s1_readdata
	wire   [1:0] mm_interconnect_0_data_a_s1_address;                         // mm_interconnect_0:data_A_s1_address -> data_A:address
	wire         mm_interconnect_0_data_a_s1_write;                           // mm_interconnect_0:data_A_s1_write -> data_A:write_n
	wire  [31:0] mm_interconnect_0_data_a_s1_writedata;                       // mm_interconnect_0:data_A_s1_writedata -> data_A:writedata
	wire         mm_interconnect_0_data_b_s1_chipselect;                      // mm_interconnect_0:data_B_s1_chipselect -> data_B:chipselect
	wire  [31:0] mm_interconnect_0_data_b_s1_readdata;                        // data_B:readdata -> mm_interconnect_0:data_B_s1_readdata
	wire   [1:0] mm_interconnect_0_data_b_s1_address;                         // mm_interconnect_0:data_B_s1_address -> data_B:address
	wire         mm_interconnect_0_data_b_s1_write;                           // mm_interconnect_0:data_B_s1_write -> data_B:write_n
	wire  [31:0] mm_interconnect_0_data_b_s1_writedata;                       // mm_interconnect_0:data_B_s1_writedata -> data_B:writedata
	wire         mm_interconnect_0_reset_pulsecounter_s1_chipselect;          // mm_interconnect_0:reset_pulseCounter_s1_chipselect -> reset_pulseCounter:chipselect
	wire  [31:0] mm_interconnect_0_reset_pulsecounter_s1_readdata;            // reset_pulseCounter:readdata -> mm_interconnect_0:reset_pulseCounter_s1_readdata
	wire   [1:0] mm_interconnect_0_reset_pulsecounter_s1_address;             // mm_interconnect_0:reset_pulseCounter_s1_address -> reset_pulseCounter:address
	wire         mm_interconnect_0_reset_pulsecounter_s1_write;               // mm_interconnect_0:reset_pulseCounter_s1_write -> reset_pulseCounter:write_n
	wire  [31:0] mm_interconnect_0_reset_pulsecounter_s1_writedata;           // mm_interconnect_0:reset_pulseCounter_s1_writedata -> reset_pulseCounter:writedata
	wire         mm_interconnect_0_wrreg_s1_chipselect;                       // mm_interconnect_0:wrreg_s1_chipselect -> wrreg:chipselect
	wire  [31:0] mm_interconnect_0_wrreg_s1_readdata;                         // wrreg:readdata -> mm_interconnect_0:wrreg_s1_readdata
	wire   [1:0] mm_interconnect_0_wrreg_s1_address;                          // mm_interconnect_0:wrreg_s1_address -> wrreg:address
	wire         mm_interconnect_0_wrreg_s1_write;                            // mm_interconnect_0:wrreg_s1_write -> wrreg:write_n
	wire  [31:0] mm_interconnect_0_wrreg_s1_writedata;                        // mm_interconnect_0:wrreg_s1_writedata -> wrreg:writedata
	wire  [31:0] mm_interconnect_0_wrfull_s1_readdata;                        // wrfull:readdata -> mm_interconnect_0:wrfull_s1_readdata
	wire   [1:0] mm_interconnect_0_wrfull_s1_address;                         // mm_interconnect_0:wrfull_s1_address -> wrfull:address
	wire  [31:0] mm_interconnect_0_screen_s1_readdata;                        // screen:readdata -> mm_interconnect_0:screen_s1_readdata
	wire   [1:0] mm_interconnect_0_screen_s1_address;                         // mm_interconnect_0:screen_s1_address -> screen:address
	wire  [31:0] mm_interconnect_0_direction_analogic_s1_readdata;            // Direction_Analogic:readdata -> mm_interconnect_0:Direction_Analogic_s1_readdata
	wire   [1:0] mm_interconnect_0_direction_analogic_s1_address;             // mm_interconnect_0:Direction_Analogic_s1_address -> Direction_Analogic:address
	wire  [31:0] mm_interconnect_0_a_s1_readdata;                             // A:readdata -> mm_interconnect_0:A_s1_readdata
	wire   [1:0] mm_interconnect_0_a_s1_address;                              // mm_interconnect_0:A_s1_address -> A:address
	wire  [31:0] mm_interconnect_0_tr_s1_readdata;                            // TR:readdata -> mm_interconnect_0:TR_s1_readdata
	wire   [1:0] mm_interconnect_0_tr_s1_address;                             // mm_interconnect_0:TR_s1_address -> TR:address
	wire  [31:0] mm_interconnect_0_tl_s1_readdata;                            // TL:readdata -> mm_interconnect_0:TL_s1_readdata
	wire   [1:0] mm_interconnect_0_tl_s1_address;                             // mm_interconnect_0:TL_s1_address -> TL:address
	wire  [31:0] mm_interconnect_0_b_s1_readdata;                             // B:readdata -> mm_interconnect_0:B_s1_readdata
	wire   [1:0] mm_interconnect_0_b_s1_address;                              // mm_interconnect_0:B_s1_address -> B:address
	wire  [31:0] mm_interconnect_0_y_s1_readdata;                             // y:readdata -> mm_interconnect_0:y_s1_readdata
	wire   [1:0] mm_interconnect_0_y_s1_address;                              // mm_interconnect_0:y_s1_address -> y:address
	wire  [31:0] mm_interconnect_0_x_s1_readdata;                             // X:readdata -> mm_interconnect_0:X_s1_readdata
	wire   [1:0] mm_interconnect_0_x_s1_address;                              // mm_interconnect_0:X_s1_address -> X:address
	wire  [31:0] mm_interconnect_0_start_s1_readdata;                         // start:readdata -> mm_interconnect_0:start_s1_readdata
	wire   [1:0] mm_interconnect_0_start_s1_address;                          // mm_interconnect_0:start_s1_address -> start:address
	wire  [31:0] mm_interconnect_0_select_button_s1_readdata;                 // select_button:readdata -> mm_interconnect_0:select_button_s1_readdata
	wire   [1:0] mm_interconnect_0_select_button_s1_address;                  // mm_interconnect_0:select_button_s1_address -> select_button:address
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [A:reset_n, B:reset_n, Direction_Analogic:reset_n, TL:reset_n, TR:reset_n, X:reset_n, data_A:reset_n, data_B:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, reset_pulseCounter:reset_n, rst_translator:in_reset, screen:reset_n, select_button:reset_n, start:reset_n, sysid_qsys_0:reset_n, wrfull:reset_n, wrreg:reset_n, y:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> rst_controller:reset_in1

	Arquitetura_A a (
		.clk      (clk_clk),                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_a_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_a_s1_readdata), //                    .readdata
		.in_port  (a_button_export)                  // external_connection.export
	);

	Arquitetura_A b (
		.clk      (clk_clk),                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_b_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_b_s1_readdata), //                    .readdata
		.in_port  (b_button_export)                  // external_connection.export
	);

	Arquitetura_Direction_Analogic direction_analogic (
		.clk      (clk_clk),                                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address  (mm_interconnect_0_direction_analogic_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_direction_analogic_s1_readdata), //                    .readdata
		.in_port  (direction_analogic_export)                         // external_connection.export
	);

	Arquitetura_A tl (
		.clk      (clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_tl_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_tl_s1_readdata), //                    .readdata
		.in_port  (tl_button_export)                  // external_connection.export
	);

	Arquitetura_A tr (
		.clk      (clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_tr_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_tr_s1_readdata), //                    .readdata
		.in_port  (tr_button_export)                  // external_connection.export
	);

	Arquitetura_A x (
		.clk      (clk_clk),                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_x_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_x_s1_readdata), //                    .readdata
		.in_port  (x_button_export)                  // external_connection.export
	);

	Arquitetura_data_A data_a (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_data_a_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_data_a_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_data_a_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_data_a_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_data_a_s1_readdata),   //                    .readdata
		.out_port   (data_a_export)                           // external_connection.export
	);

	Arquitetura_data_A data_b (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_data_b_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_data_b_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_data_b_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_data_b_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_data_b_s1_readdata),   //                    .readdata
		.out_port   (data_b_export)                           // external_connection.export
	);

	Arquitetura_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	Arquitetura_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	Arquitetura_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	Arquitetura_reset_pulseCounter reset_pulsecounter (
		.clk        (clk_clk),                                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_reset_pulsecounter_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reset_pulsecounter_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reset_pulsecounter_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reset_pulsecounter_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reset_pulsecounter_s1_readdata),   //                    .readdata
		.out_port   (reset_pulsecounter_export)                           // external_connection.export
	);

	Arquitetura_A screen (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_screen_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_screen_s1_readdata), //                    .readdata
		.in_port  (screen_export)                         // external_connection.export
	);

	Arquitetura_A select_button (
		.clk      (clk_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_select_button_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_select_button_s1_readdata), //                    .readdata
		.in_port  (select_button_export)                         // external_connection.export
	);

	Arquitetura_A start (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_start_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_start_s1_readdata), //                    .readdata
		.in_port  (start_button_export)                  // external_connection.export
	);

	Arquitetura_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	Arquitetura_A wrfull (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_wrfull_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_wrfull_s1_readdata), //                    .readdata
		.in_port  (wrfull_export)                         // external_connection.export
	);

	Arquitetura_reset_pulseCounter wrreg (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_wrreg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_wrreg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_wrreg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_wrreg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_wrreg_s1_readdata),   //                    .readdata
		.out_port   (wrreg_export)                           // external_connection.export
	);

	Arquitetura_A y (
		.clk      (clk_clk),                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_y_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_y_s1_readdata), //                    .readdata
		.in_port  (y_button_export)                  // external_connection.export
	);

	Arquitetura_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.A_s1_address                                   (mm_interconnect_0_a_s1_address),                              //                                     A_s1.address
		.A_s1_readdata                                  (mm_interconnect_0_a_s1_readdata),                             //                                         .readdata
		.B_s1_address                                   (mm_interconnect_0_b_s1_address),                              //                                     B_s1.address
		.B_s1_readdata                                  (mm_interconnect_0_b_s1_readdata),                             //                                         .readdata
		.data_A_s1_address                              (mm_interconnect_0_data_a_s1_address),                         //                                data_A_s1.address
		.data_A_s1_write                                (mm_interconnect_0_data_a_s1_write),                           //                                         .write
		.data_A_s1_readdata                             (mm_interconnect_0_data_a_s1_readdata),                        //                                         .readdata
		.data_A_s1_writedata                            (mm_interconnect_0_data_a_s1_writedata),                       //                                         .writedata
		.data_A_s1_chipselect                           (mm_interconnect_0_data_a_s1_chipselect),                      //                                         .chipselect
		.data_B_s1_address                              (mm_interconnect_0_data_b_s1_address),                         //                                data_B_s1.address
		.data_B_s1_write                                (mm_interconnect_0_data_b_s1_write),                           //                                         .write
		.data_B_s1_readdata                             (mm_interconnect_0_data_b_s1_readdata),                        //                                         .readdata
		.data_B_s1_writedata                            (mm_interconnect_0_data_b_s1_writedata),                       //                                         .writedata
		.data_B_s1_chipselect                           (mm_interconnect_0_data_b_s1_chipselect),                      //                                         .chipselect
		.Direction_Analogic_s1_address                  (mm_interconnect_0_direction_analogic_s1_address),             //                    Direction_Analogic_s1.address
		.Direction_Analogic_s1_readdata                 (mm_interconnect_0_direction_analogic_s1_readdata),            //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.reset_pulseCounter_s1_address                  (mm_interconnect_0_reset_pulsecounter_s1_address),             //                    reset_pulseCounter_s1.address
		.reset_pulseCounter_s1_write                    (mm_interconnect_0_reset_pulsecounter_s1_write),               //                                         .write
		.reset_pulseCounter_s1_readdata                 (mm_interconnect_0_reset_pulsecounter_s1_readdata),            //                                         .readdata
		.reset_pulseCounter_s1_writedata                (mm_interconnect_0_reset_pulsecounter_s1_writedata),           //                                         .writedata
		.reset_pulseCounter_s1_chipselect               (mm_interconnect_0_reset_pulsecounter_s1_chipselect),          //                                         .chipselect
		.screen_s1_address                              (mm_interconnect_0_screen_s1_address),                         //                                screen_s1.address
		.screen_s1_readdata                             (mm_interconnect_0_screen_s1_readdata),                        //                                         .readdata
		.select_button_s1_address                       (mm_interconnect_0_select_button_s1_address),                  //                         select_button_s1.address
		.select_button_s1_readdata                      (mm_interconnect_0_select_button_s1_readdata),                 //                                         .readdata
		.start_s1_address                               (mm_interconnect_0_start_s1_address),                          //                                 start_s1.address
		.start_s1_readdata                              (mm_interconnect_0_start_s1_readdata),                         //                                         .readdata
		.sysid_qsys_0_control_slave_address             (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),       //                                         .readdata
		.TL_s1_address                                  (mm_interconnect_0_tl_s1_address),                             //                                    TL_s1.address
		.TL_s1_readdata                                 (mm_interconnect_0_tl_s1_readdata),                            //                                         .readdata
		.TR_s1_address                                  (mm_interconnect_0_tr_s1_address),                             //                                    TR_s1.address
		.TR_s1_readdata                                 (mm_interconnect_0_tr_s1_readdata),                            //                                         .readdata
		.wrfull_s1_address                              (mm_interconnect_0_wrfull_s1_address),                         //                                wrfull_s1.address
		.wrfull_s1_readdata                             (mm_interconnect_0_wrfull_s1_readdata),                        //                                         .readdata
		.wrreg_s1_address                               (mm_interconnect_0_wrreg_s1_address),                          //                                 wrreg_s1.address
		.wrreg_s1_write                                 (mm_interconnect_0_wrreg_s1_write),                            //                                         .write
		.wrreg_s1_readdata                              (mm_interconnect_0_wrreg_s1_readdata),                         //                                         .readdata
		.wrreg_s1_writedata                             (mm_interconnect_0_wrreg_s1_writedata),                        //                                         .writedata
		.wrreg_s1_chipselect                            (mm_interconnect_0_wrreg_s1_chipselect),                       //                                         .chipselect
		.X_s1_address                                   (mm_interconnect_0_x_s1_address),                              //                                     X_s1.address
		.X_s1_readdata                                  (mm_interconnect_0_x_s1_readdata),                             //                                         .readdata
		.y_s1_address                                   (mm_interconnect_0_y_s1_address),                              //                                     y_s1.address
		.y_s1_readdata                                  (mm_interconnect_0_y_s1_readdata)                              //                                         .readdata
	);

	Arquitetura_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
